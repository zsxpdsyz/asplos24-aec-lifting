`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  wire [0:0] PI_clk = clock;
  cva6_lsu_formal UUT (
    .clk(PI_clk)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$formal$cva6_lsu_formal.\v:173$10_EN  = 1'b0;
    // UUT.$formal$cva6_lsu_formal.\v:210$12_CHECK  = 1'b0;
    UUT.counter = 3'b000;
    UUT.init = 1'b1;
    UUT.local_ready_1 = 1'b0;
    UUT.local_ready_2 = 1'b0;
    UUT.pc_1 = 32'b00000000000000000000000000000000;
    UUT.pc_2 = 32'b00000000000000000000000000000000;
    UUT.reset = 1'b1;
    UUT.shim_i_1.load_cooldown = 3'b000;
    UUT.shim_i_1.loadstore_addr = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.loadstore_fsm = 3'b000;
    UUT.shim_i_1.loadstore_state = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10690  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10692  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10694  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10696  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10698  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10700  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10702  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10704  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10706  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10708  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10710  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10712  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10714  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10716  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10718  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10720  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10722  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10724  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10726  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10728  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10730  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10732  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10734  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10736  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10738  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10740  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10742  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10744  = 2'b00;
    UUT.shim_i_1.\mem[0]  = 32'b11111111111111111111001111100011;
    UUT.shim_i_1.\mem[10]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[11]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[12]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[13]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[14]  = 32'b11111111111111111111100001000111;
    UUT.shim_i_1.\mem[15]  = 32'b11111111111111111111000100111011;
    UUT.shim_i_1.\mem[16]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[18]  = 32'b11111111111111111111011011101111;
    UUT.shim_i_1.\mem[19]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[1]  = 32'b11111111111111111111010110111111;
    UUT.shim_i_1.\mem[20]  = 32'b11111111111111111111111111101111;
    UUT.shim_i_1.\mem[21]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[22]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[23]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[24]  = 32'b11111111111111111111011011101111;
    UUT.shim_i_1.\mem[25]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[26]  = 32'b11111111111111111111010010001110;
    UUT.shim_i_1.\mem[27]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[28]  = 32'b11111111111111111111000010111111;
    UUT.shim_i_1.\mem[29]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[2]  = 32'b11111111111111111111111110011001;
    UUT.shim_i_1.\mem[30]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[31]  = 32'b11111111111111111111110001110111;
    UUT.shim_i_1.\mem[3]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[4]  = 32'b11111111111111111111000010111111;
    UUT.shim_i_1.\mem[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[6]  = 32'b11111111111111111111101111011001;
    UUT.shim_i_1.\mem[7]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[8]  = 32'b11111111111111111111001010111111;
    UUT.shim_i_1.\mem[9]  = 32'b11111111111111111110001010111111;
    UUT.shim_i_1.ready_o = 1'b0;
    UUT.shim_i_1.\regfile[0]  = 32'b01111111111111111111010010111111;
    UUT.shim_i_1.\regfile[10]  = 32'b11111111111111111111100101101000;
    UUT.shim_i_1.\regfile[11]  = 32'b11111111111111111111011001110110;
    UUT.shim_i_1.\regfile[12]  = 32'b11111111111111111111011000001100;
    UUT.shim_i_1.\regfile[13]  = 32'b11111111111111111111010101010000;
    UUT.shim_i_1.\regfile[14]  = 32'b11111111111111111110111110000001;
    UUT.shim_i_1.\regfile[15]  = 32'b11111111111111111111101010100001;
    UUT.shim_i_1.\regfile[16]  = 32'b11111111111111111111010010001110;
    UUT.shim_i_1.\regfile[17]  = 32'b11111111111111111110101001100100;
    UUT.shim_i_1.\regfile[18]  = 32'b11111111111111111111010010111111;
    UUT.shim_i_1.\regfile[19]  = 32'b11111111111111111111001100000101;
    UUT.shim_i_1.\regfile[1]  = 32'b11111111111111111110110100101011;
    UUT.shim_i_1.\regfile[20]  = 32'b01111111111111111110110100111010;
    UUT.shim_i_1.\regfile[21]  = 32'b01111111111111111110001010001000;
    UUT.shim_i_1.\regfile[22]  = 32'b01111111111111111110110111111001;
    UUT.shim_i_1.\regfile[23]  = 32'b11111111111111111111111000011011;
    UUT.shim_i_1.\regfile[24]  = 32'b10000000000000000000000000101000;
    UUT.shim_i_1.\regfile[25]  = 32'b11111111111111111111101000011010;
    UUT.shim_i_1.\regfile[26]  = 32'b01111111111111111110111000011000;
    UUT.shim_i_1.\regfile[27]  = 32'b11111111111111111111100010011010;
    UUT.shim_i_1.\regfile[28]  = 32'b11111111111111111111001100000010;
    UUT.shim_i_1.\regfile[29]  = 32'b11111111111111111111111100001001;
    UUT.shim_i_1.\regfile[2]  = 32'b01111111111111111110111110101110;
    UUT.shim_i_1.\regfile[30]  = 32'b11111111111111111110000010111001;
    UUT.shim_i_1.\regfile[31]  = 32'b11111111111111111110110000001001;
    UUT.shim_i_1.\regfile[3]  = 32'b11111111111111111111010110111011;
    UUT.shim_i_1.\regfile[4]  = 32'b11111111111111111111001110111101;
    UUT.shim_i_1.\regfile[5]  = 32'b11111111111111111111011111100000;
    UUT.shim_i_1.\regfile[6]  = 32'b11111111111111111111001100010100;
    UUT.shim_i_1.\regfile[7]  = 32'b11111111111111111110100000001000;
    UUT.shim_i_1.\regfile[8]  = 32'b11111111111111111111011100011010;
    UUT.shim_i_1.\regfile[9]  = 32'b11111111111111111111111101101000;
    UUT.shim_i_1.store_cooldown = 1'b0;
    UUT.shim_i_1.store_count = 3'b000;
    UUT.shim_i_1.store_uncommitted = 1'b0;
    UUT.shim_i_1.tb_io_instr_i = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.tb_io_instr_valid_i = 1'b0;
    UUT.shim_i_1.tb_io_is_load_i = 1'b0;
    UUT.shim_i_1.tb_io_load_mem_resp_i = 1'b0;
    UUT.shim_i_1.tb_io_store_commit_i = 1'b0;
    UUT.shim_i_1.tb_io_store_mem_resp_i = 1'b0;
    UUT.shim_i_2.load_cooldown = 3'b000;
    UUT.shim_i_2.loadstore_addr = 32'b00000000000000000000000000000000;
    UUT.shim_i_2.loadstore_fsm = 3'b000;
    UUT.shim_i_2.loadstore_state = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10690  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10692  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10694  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10696  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10698  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10700  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10702  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10704  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10706  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10708  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10710  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10712  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10714  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10716  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10718  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10720  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10722  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10724  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10726  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10728  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10730  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10732  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10734  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10736  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10738  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10740  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10742  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10744  = 2'b00;
    UUT.shim_i_2.\mem[0]  = 32'b11111111111111111111001111100011;
    UUT.shim_i_2.\mem[10]  = 32'b11111111111111111111111101101000;
    UUT.shim_i_2.\mem[11]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[12]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[13]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[14]  = 32'b11111111111111111110101111111111;
    UUT.shim_i_2.\mem[15]  = 32'b11111111111111111111011100101101;
    UUT.shim_i_2.\mem[16]  = 32'b11111111111111111111010101101011;
    UUT.shim_i_2.\mem[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[18]  = 32'b11111111111111111111001101001001;
    UUT.shim_i_2.\mem[19]  = 32'b11111111111111111111110011111011;
    UUT.shim_i_2.\mem[1]  = 32'b11111111111111111111000110111011;
    UUT.shim_i_2.\mem[20]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[21]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[22]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[23]  = 32'b11111111111111111111011010111111;
    UUT.shim_i_2.\mem[24]  = 32'b11111111111111111111001101001001;
    UUT.shim_i_2.\mem[25]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[26]  = 32'b11111111111111111111111111001011;
    UUT.shim_i_2.\mem[27]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[28]  = 32'b11111111111111111111100010000010;
    UUT.shim_i_2.\mem[29]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[2]  = 32'b11111111111111111111111111101011;
    UUT.shim_i_2.\mem[30]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[31]  = 32'b11111111111111111111110001110111;
    UUT.shim_i_2.\mem[3]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[4]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[6]  = 32'b11111111111111111111011111101101;
    UUT.shim_i_2.\mem[7]  = 32'b11111111111111111111111110011001;
    UUT.shim_i_2.\mem[8]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[9]  = 32'b11111111111111111110101101000011;
    UUT.shim_i_2.ready_o = 1'b0;
    UUT.shim_i_2.\regfile[0]  = 32'b01111111111111111111010010111111;
    UUT.shim_i_2.\regfile[10]  = 32'b11111111111111111111100101101000;
    UUT.shim_i_2.\regfile[11]  = 32'b11111111111111111111011001110110;
    UUT.shim_i_2.\regfile[12]  = 32'b11111111111111111111011000001100;
    UUT.shim_i_2.\regfile[13]  = 32'b11111111111111111111010101010000;
    UUT.shim_i_2.\regfile[14]  = 32'b11111111111111111110111110000001;
    UUT.shim_i_2.\regfile[15]  = 32'b11111111111111111111101010100001;
    UUT.shim_i_2.\regfile[16]  = 32'b11111111111111111111010010001110;
    UUT.shim_i_2.\regfile[17]  = 32'b11111111111111111110101001100100;
    UUT.shim_i_2.\regfile[18]  = 32'b11111111111111111111010010111111;
    UUT.shim_i_2.\regfile[19]  = 32'b11111111111111111111001100000101;
    UUT.shim_i_2.\regfile[1]  = 32'b11111111111111111110110100101011;
    UUT.shim_i_2.\regfile[20]  = 32'b01111111111111111110110100111010;
    UUT.shim_i_2.\regfile[21]  = 32'b01111111111111111110001010001000;
    UUT.shim_i_2.\regfile[22]  = 32'b01111111111111111110110111111001;
    UUT.shim_i_2.\regfile[23]  = 32'b11111111111111111111111000011011;
    UUT.shim_i_2.\regfile[24]  = 32'b10000000000000000000000000101000;
    UUT.shim_i_2.\regfile[25]  = 32'b11111111111111111111101000011010;
    UUT.shim_i_2.\regfile[26]  = 32'b01111111111111111110111000011000;
    UUT.shim_i_2.\regfile[27]  = 32'b11111111111111111111100010011010;
    UUT.shim_i_2.\regfile[28]  = 32'b11111111111111111111001100000010;
    UUT.shim_i_2.\regfile[29]  = 32'b11111111111111111111111100001001;
    UUT.shim_i_2.\regfile[2]  = 32'b01111111111111111110111110101110;
    UUT.shim_i_2.\regfile[30]  = 32'b11111111111111111110000010111001;
    UUT.shim_i_2.\regfile[31]  = 32'b11111111111111111110110000001001;
    UUT.shim_i_2.\regfile[3]  = 32'b11111111111111111111010110111011;
    UUT.shim_i_2.\regfile[4]  = 32'b11111111111111111111001110111101;
    UUT.shim_i_2.\regfile[5]  = 32'b11111111111111111111011111100000;
    UUT.shim_i_2.\regfile[6]  = 32'b11111111111111111111001100010100;
    UUT.shim_i_2.\regfile[7]  = 32'b11111111111111111110100000001000;
    UUT.shim_i_2.\regfile[8]  = 32'b11111111111111111111011100011010;
    UUT.shim_i_2.\regfile[9]  = 32'b11111111111111111111111101101000;
    UUT.shim_i_2.store_cooldown = 1'b0;
    UUT.shim_i_2.store_count = 3'b000;
    UUT.shim_i_2.store_uncommitted = 1'b0;
    UUT.shim_i_2.tb_io_instr_i = 32'b00000000000000000000000000000000;
    UUT.shim_i_2.tb_io_instr_valid_i = 1'b0;
    UUT.shim_i_2.tb_io_is_load_i = 1'b0;
    UUT.shim_i_2.tb_io_load_mem_resp_i = 1'b0;
    UUT.shim_i_2.tb_io_store_commit_i = 1'b0;
    UUT.shim_i_2.tb_io_store_mem_resp_i = 1'b0;
    UUT.tb_io_instr_i_1 = 32'b01100100000011000000100000000011;
    UUT.tb_io_instr_i_2 = 32'b00000001000011001001010010000011;
    UUT.tb_io_instr_valid_i_1 = 1'b1;
    UUT.tb_io_instr_valid_i_2 = 1'b1;
    UUT.instr2 = 32'b00011100011111010010111110000011;
    UUT.instr1 = 32'b11110010000000000010111010100011;
    UUT.instr0 = 32'b11110100111011110010000110000011;
    UUT.instr3 = 32'b11010011110011111010000000000011;

    // state 0
    UUT.tb_io_store_mem_resp_i_2 = 1'b0;
    UUT.tb_io_store_mem_resp_i_1 = 1'b0;
    UUT.tb_io_load_mem_resp_i_2 = 1'b0;
    UUT.tb_io_load_mem_resp_i_1 = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 4
    if (cycle == 3) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 5
    if (cycle == 4) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 6
    if (cycle == 5) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 7
    if (cycle == 6) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 8
    if (cycle == 7) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 9
    if (cycle == 8) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 10
    if (cycle == 9) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 11
    if (cycle == 10) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 12
    if (cycle == 11) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 13
    if (cycle == 12) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 14
    if (cycle == 13) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 15
    if (cycle == 14) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 16
    if (cycle == 15) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 17
    if (cycle == 16) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 18
    if (cycle == 17) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 19
    if (cycle == 18) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 20
    if (cycle == 19) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 21
    if (cycle == 20) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 22
    if (cycle == 21) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 23
    if (cycle == 22) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 24
    if (cycle == 23) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 25
    if (cycle == 24) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 26
    if (cycle == 25) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 27
    if (cycle == 26) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 28
    if (cycle == 27) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 29
    if (cycle == 28) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 30
    if (cycle == 29) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 31
    if (cycle == 30) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 32
    if (cycle == 31) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 33
    if (cycle == 32) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 34
    if (cycle == 33) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 35
    if (cycle == 34) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 36
    if (cycle == 35) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 37
    if (cycle == 36) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 38
    if (cycle == 37) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    genclock <= cycle < 38;
    cycle <= cycle + 1;
  end
endmodule
