`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  wire [0:0] PI_clk = clock;
  cva6_lsu_formal UUT (
    .clk(PI_clk)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$formal$cva6_lsu_formal.\v:169$7_EN  = 1'b0;
    // UUT.$formal$cva6_lsu_formal.\v:206$9_CHECK  = 1'b0;
    UUT.counter = 3'b000;
    UUT.init = 1'b1;
    UUT.local_ready_1 = 1'b0;
    UUT.local_ready_2 = 1'b0;
    UUT.pc_1 = 32'b00000000000000000000000000000000;
    UUT.pc_2 = 32'b00000000000000000000000000000000;
    UUT.reset = 1'b1;
    UUT.shim_i_1.load_cooldown = 3'b000;
    UUT.shim_i_1.loadstore_addr = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.loadstore_fsm = 3'b000;
    UUT.shim_i_1.loadstore_state = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10645  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10647  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10649  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10651  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10653  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10655  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10657  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10659  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10661  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10663  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10665  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10667  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10669  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10671  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10673  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10675  = 1'b0;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10677  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10679  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10681  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10683  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10685  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10687  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10689  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10691  = 8'b00000000;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10693  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10695  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10697  = 2'b00;
    // UUT.shim_i_1.lsu_model_i.$auto$async2sync.\cc:140:execute$10699  = 2'b00;
    UUT.shim_i_1.\mem[0]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[10]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[11]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[12]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[13]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[14]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[15]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[16]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[18]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[19]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[1]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[20]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[21]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[22]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[23]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[24]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[25]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[26]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[27]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[28]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[29]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[2]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[30]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[31]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[3]  = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.\mem[4]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[6]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[7]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[8]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\mem[9]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.ready_o = 1'b0;
    UUT.shim_i_1.\regfile[0]  = 32'b00111111111111111111110011101000;
    UUT.shim_i_1.\regfile[10]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[11]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[12]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[13]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[14]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[15]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[16]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[18]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[19]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[1]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[20]  = 32'b11111111111111111111101111001011;
    UUT.shim_i_1.\regfile[21]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[22]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[23]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[24]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[25]  = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.\regfile[26]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[27]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[28]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[29]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[2]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[30]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[31]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[3]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[4]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[6]  = 32'b11111111111111111111010100000111;
    UUT.shim_i_1.\regfile[7]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[8]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.\regfile[9]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_1.store_cooldown = 1'b0;
    UUT.shim_i_1.store_count = 3'b000;
    UUT.shim_i_1.store_uncommitted = 1'b0;
    UUT.shim_i_1.tb_io_instr_i = 32'b00000000000000000000000000000000;
    UUT.shim_i_1.tb_io_instr_valid_i = 1'b0;
    UUT.shim_i_1.tb_io_is_load_i = 1'b0;
    UUT.shim_i_1.tb_io_load_mem_resp_i = 1'b0;
    UUT.shim_i_1.tb_io_store_commit_i = 1'b0;
    UUT.shim_i_1.tb_io_store_mem_resp_i = 1'b0;
    UUT.shim_i_2.load_cooldown = 3'b000;
    UUT.shim_i_2.loadstore_addr = 32'b00000000000000000000000000000000;
    UUT.shim_i_2.loadstore_fsm = 3'b000;
    UUT.shim_i_2.loadstore_state = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10645  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10647  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10649  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10651  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10653  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10655  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10657  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10659  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10661  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10663  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10665  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10667  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10669  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10671  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10673  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10675  = 1'b0;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10677  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10679  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10681  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10683  = 32'b00000000000000000000000000000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10685  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10687  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10689  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10691  = 8'b00000000;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10693  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10695  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10697  = 2'b00;
    // UUT.shim_i_2.lsu_model_i.$auto$async2sync.\cc:140:execute$10699  = 2'b00;
    UUT.shim_i_2.\mem[0]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[10]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[11]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[12]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[13]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[14]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[15]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[16]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[18]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[19]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[1]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[20]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[21]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[22]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[23]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[24]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[25]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[26]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[27]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[28]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[29]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[2]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[30]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[31]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[3]  = 32'b00000000000000000000000000000000;
    UUT.shim_i_2.\mem[4]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[6]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[7]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[8]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\mem[9]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.ready_o = 1'b0;
    UUT.shim_i_2.\regfile[0]  = 32'b11111111111111111110110011100100;
    UUT.shim_i_2.\regfile[10]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[11]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[12]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[13]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[14]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[15]  = 32'b01111111111111111111111111111111;
    UUT.shim_i_2.\regfile[16]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[17]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[18]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[19]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[1]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[20]  = 32'b11111111111111111111010001001011;
    UUT.shim_i_2.\regfile[21]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[22]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[23]  = 32'b10000000000000000000000000000000;
    UUT.shim_i_2.\regfile[24]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[25]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[26]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[27]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[28]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[29]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[2]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[30]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[31]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[3]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[4]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[5]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[6]  = 32'b10000000000000000000010011111111;
    UUT.shim_i_2.\regfile[7]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[8]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.\regfile[9]  = 32'b11111111111111111111111111111111;
    UUT.shim_i_2.store_cooldown = 1'b0;
    UUT.shim_i_2.store_count = 3'b000;
    UUT.shim_i_2.store_uncommitted = 1'b0;
    UUT.shim_i_2.tb_io_instr_i = 32'b00000000000000000000000000000000;
    UUT.shim_i_2.tb_io_instr_valid_i = 1'b0;
    UUT.shim_i_2.tb_io_is_load_i = 1'b0;
    UUT.shim_i_2.tb_io_load_mem_resp_i = 1'b0;
    UUT.shim_i_2.tb_io_store_commit_i = 1'b0;
    UUT.shim_i_2.tb_io_store_mem_resp_i = 1'b0;
    UUT.tb_io_instr_i_1 = 32'b01000000000000000100110010010011;
    UUT.tb_io_instr_i_2 = 32'b01000100000110110100101110010011;
    UUT.tb_io_instr_valid_i_1 = 1'b0;
    UUT.tb_io_instr_valid_i_2 = 1'b0;
    UUT.instr2 = 32'b10110000000000110010000000000011;
    UUT.instr1 = 32'b00110000000000000010111000100011;
    UUT.instr0 = 32'b11000100001110100010010010000011;
    UUT.instr3 = 32'b00000000000000000000000000010011;

    // state 0
    UUT.tb_io_store_mem_resp_i_2 = 1'b0;
    UUT.tb_io_store_mem_resp_i_1 = 1'b0;
    UUT.tb_io_load_mem_resp_i_2 = 1'b0;
    UUT.tb_io_load_mem_resp_i_1 = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 4
    if (cycle == 3) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 5
    if (cycle == 4) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 6
    if (cycle == 5) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 7
    if (cycle == 6) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 8
    if (cycle == 7) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 9
    if (cycle == 8) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 10
    if (cycle == 9) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 11
    if (cycle == 10) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 12
    if (cycle == 11) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 13
    if (cycle == 12) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 14
    if (cycle == 13) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 15
    if (cycle == 14) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 16
    if (cycle == 15) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 17
    if (cycle == 16) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 18
    if (cycle == 17) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 19
    if (cycle == 18) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 20
    if (cycle == 19) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 21
    if (cycle == 20) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 22
    if (cycle == 21) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 23
    if (cycle == 22) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 24
    if (cycle == 23) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 25
    if (cycle == 24) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 26
    if (cycle == 25) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 27
    if (cycle == 26) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 28
    if (cycle == 27) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    // state 29
    if (cycle == 28) begin
      UUT.tb_io_store_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_store_mem_resp_i_1 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_2 <= 1'b0;
      UUT.tb_io_load_mem_resp_i_1 <= 1'b0;
    end

    genclock <= cycle < 29;
    cycle <= cycle + 1;
  end
endmodule
